`ifdef FIBONACCI
    `define BENCHMARK "fibonacci_p.v"
`else
    `define BENCHMARK "test_instr.txt"
`endif

